module hello;
 initial begin
    $display("Helllo Verilog!");
 end 
endmodule